
module vga_char_86x32 #(
    parameter VGA_CLK_DIV = 1
)(
    // clock and reset
	input  logic         clk, rst_n,
    // vga interfaces
	output logic         hsync, vsync,
	output logic         red, green, blue,
    // ascii read interface
    output logic         req,
    output logic [ 6:0]  reqx,
    output logic [ 4:0]  reqy,
    input  logic [ 6:0]  ascii
);

localparam  H_END           =                 10'd688,
            H_BRSTART       = H_END         + 10'd4  ,
            H_BREND         = H_BRSTART     + 10'd30 ,
            H_SYNCSTART     = H_BREND       + 10'd25 ,
            H_SYNCEND       = H_SYNCSTART   + 10'd128,
            H_BLSTART       = H_SYNCEND     + 10'd89 ,
            H_BLEND         = H_BLSTART     + 10'd30 ,
            H_PERIOD        = H_BLEND       + 10'd4  ,
            V_END           =                 10'd512,
            V_BRSTART       = V_END         + 10'd4  ,
            V_BREND         = V_BRSTART     + 10'd30 ,
            V_SYNCSTART     = V_BREND       + 10'd38 ,
            V_SYNCEND       = V_SYNCSTART   + 10'd4  ,
            V_BLSTART       = V_SYNCEND     + 10'd66 ,
            V_BLEND         = V_BLSTART     + 10'd30 ,
            V_PERIOD        = V_BLEND       + 10'd4  ;

logic [3:0] rlp=4'h0, clp=4'h0, hsp=4'h0, vsp=4'h0;
logic vlbr=1'b0, vgbl=1'b0, vlbl=1'b0, vgbr=1'b0, hlbr=1'b0, hgbl=1'b0, hlbl=1'b0, hgbr=1'b0;
logic vir=1'b0, hir=1'b0, vbr=1'b0, hbr=1'b0, vbl=1'b0, hbl=1'b0, hb=1'b0, vb=1'b0, border=1'b0;
logic [9:0] cnt = 0, hcnt = 0, vcnt = 0;
logic req1 = 1'b0, req2 = 1'b0;
logic [6:0] ascii_bufferout, ascii_latch=8'h0, ascii_to_rom;
logic [7:0] rom_data;
logic [6:0] x_h, x_h1=7'h0, x_h2=7'h0;
logic [5:0] y_h;

logic [2:0] x_l, x_l1 = 3'h0, x_l2 = 3'h0, x_l3 = 3'h0, x_l4 = 3'h0;
logic [3:0] y_l, y_l1 = 4'h0, y_l2 = 4'h0, y_l3 = 4'h0;

assign {x_h, x_l} = hcnt;
assign {y_h, y_l} = vcnt;

initial begin hsync=1'b0; vsync=1'b0; {red,green,blue}=3'h0; req=1'b0; {reqx, reqy} = '0; end

always @ (posedge clk)
    if(~rst_n) begin
        vlbr<= 1'b0;
        vgbl<= 1'b0;
        vlbl<= 1'b0;
        vgbr<= 1'b0;
        hlbr<= 1'b0;
        hgbl<= 1'b0;
        hlbl<= 1'b0;
        hgbr<= 1'b0;
        vir <= 1'b0;
        hir <= 1'b0;
        vbr <= 1'b0;
        hbr <= 1'b0;
        vbl <= 1'b0;
        hbl <= 1'b0;
        hb  <= 1'b0;
        vb  <= 1'b0;
        border <= 1'b0;
    end else begin
        vlbr<= vcnt <  V_BREND  ;
        vgbl<= vcnt >= V_BLSTART;
        vlbl<= vcnt <  V_BLEND  ;
        vgbr<= vcnt >= V_BRSTART;
        hlbr<= hcnt <  H_BREND  ;
        hgbl<= hcnt >= H_BLSTART;
        hlbl<= hcnt <  H_BLEND;
        hgbr<= hcnt >= H_BRSTART;
        vir <= vlbr | vgbl;
        hir <= hlbr | hgbl;
        vbr <= vgbr & vlbr;
        hbr <= hgbr & hlbr;
        vbl <= vgbl & vlbl;
        hbl <= hgbl & hlbl;
        hb  <= (hbr | hbl) & vir;
        vb  <= (vbr | vbl) & hir;
        border <= hb | vb;
    end

always @ (posedge clk or negedge rst_n)
    if(~rst_n) begin
        cnt  <= 10'h0;
        hcnt <= 10'h0;
        vcnt <= 10'h0;
    end else begin
        cnt <= (cnt<(VGA_CLK_DIV-1)) ? cnt + 10'h1 : 10'h0;
        if(cnt==10'h0) begin
            if(hcnt < H_PERIOD) begin
                hcnt <= hcnt + 10'h1;
            end else begin
                hcnt <= 10'h0;
                vcnt <= (vcnt<V_PERIOD) ? vcnt + 10'h1 : 10'h0;
            end
        end
    end
    
always @ (posedge clk or negedge rst_n)
    if(~rst_n) begin
        req <= 1'b0;
        req1<= 1'b0;
        req2<= 1'b0;
    end else begin
        req <= cnt==10'h0 && hcnt<H_END && vcnt<V_END && x_l==3'h0 && y_l==4'h0;
        req1<= req;
        req2<= req1;
    end
    
always @ (posedge clk or negedge rst_n)
    if(~rst_n) begin
        clp <= 4'h0;
        rlp <= 4'h0;
        hsp <= 4'h0;
        vsp <= 4'h0;
    end else begin
        clp <= {clp[2:0], ( cnt==10'h0 ) };
        rlp <= {rlp[2:0], ( hcnt<H_END && vcnt<V_END ) };
        hsp <= {hsp[2:0], ( hcnt>=H_SYNCSTART && hcnt<H_SYNCEND ) };
        vsp <= {vsp[2:0], ( vcnt>=V_SYNCSTART && vcnt<V_SYNCEND ) };
    end

always @ (posedge clk or negedge rst_n)
    if(~rst_n) begin
        {reqy, reqx} <= '0;
    end else begin
        if( cnt==10'h0 && hcnt<H_END && vcnt<V_END ) begin
            {reqy, reqx} <= {y_h[4:0],x_h};
        end else begin
            {reqy, reqx} <= '0;
        end
    end
    
always @ (posedge clk or negedge rst_n)
    if(~rst_n)
        {x_l1, y_l1, x_l2, y_l2, x_l3, y_l3, x_l4, x_h1, x_h2} <= 38'h0;
    else
        {x_l1, y_l1, x_l2, y_l2, x_l3, y_l3, x_l4, x_h1, x_h2} <= {x_l, y_l, x_l1, y_l1, x_l2, y_l2, x_l3, x_h, x_h1};

always @ (posedge clk or negedge rst_n)
    if(~rst_n) begin
        hsync <= 1'b0;
        vsync <= 1'b0;
        {red,green,blue} <= 3'h0;
    end else begin
        if(clp[3]) begin
            hsync <= ~hsp[3];
            vsync <= ~vsp[3];
            if(rlp[3])
                {red,green,blue} <= {3{rom_data[x_l4]}};
            else if(border)
                {red,green,blue} <= 3'b100;
            else
                {red,green,blue} <= 3'b000;
        end
    end
    
always @ (posedge clk or negedge rst_n)
    if(~rst_n)
        ascii_latch <= 6'h0;
    else begin
        ascii_latch <= req1 ? ascii : 6'h0;
    end

assign ascii_to_rom = req2 ? ascii_latch : ascii_bufferout;

// buffered a line(86 chars), The goal is to minimize the number of memory accesses
ram128B vga_line_buffer_i(            // 128B
    .clk        (  clk                 ),
    .i_we       (  req1                ),
    .i_addr     (  x_h2                ),
    .i_wdata    (  ascii               ),
    .o_rdata    (  ascii_bufferout     )
);

char8x16_rom char_8x16_rom_i(
    .clk        ( clk                  ),
    .addr       ( {ascii_to_rom, y_l3} ),
    .data       ( rom_data             )
);

endmodule













module ram128B(            // 128B
    input  logic        clk,
    input  logic        i_we,
    input  logic [ 6:0] i_addr,
    input  logic [ 6:0] i_wdata,
    output logic [ 6:0] o_rdata
);
initial o_rdata = 7'h0;

logic [6:0] data_ram_cell [0:127];
    
always @ (posedge clk)
    o_rdata <= data_ram_cell[i_addr];

always @ (posedge clk)
    if(i_we) 
        data_ram_cell[i_addr] <= i_wdata;

endmodule













module char8x16_rom(
    input  logic        clk,
    input  logic [10:0] addr,
    output logic [ 7:0] data
);

wire [0:2047] [7:0] rom_cell = {
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h18,
    8'h18,
    8'h18,
    8'h18,
    8'h18,
    8'h18,
    8'h10,
    8'h00,
    8'h10,
    8'h18,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h2c,
    8'h24,
    8'h24,
    8'h24,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h68,
    8'h24,
    8'hfe,
    8'h24,
    8'h24,
    8'h24,
    8'h7e,
    8'h24,
    8'h24,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h10,
    8'h7c,
    8'h16,
    8'h12,
    8'h16,
    8'h38,
    8'h68,
    8'h48,
    8'h48,
    8'h3e,
    8'h08,
    8'h08,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h86,
    8'h4b,
    8'h69,
    8'h2e,
    8'h10,
    8'h08,
    8'h68,
    8'h94,
    8'h92,
    8'h63,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h3c,
    8'h26,
    8'h26,
    8'h1c,
    8'h4e,
    8'h52,
    8'h73,
    8'h62,
    8'hfe,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h18,
    8'h18,
    8'h18,
    8'h18,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h20,
    8'h10,
    8'h18,
    8'h08,
    8'h0c,
    8'h0c,
    8'h0c,
    8'h0c,
    8'h08,
    8'h08,
    8'h18,
    8'h30,
    8'h20,
    8'h00,
    8'h00,
    8'h00,
    8'h04,
    8'h08,
    8'h10,
    8'h10,
    8'h30,
    8'h20,
    8'h20,
    8'h20,
    8'h30,
    8'h10,
    8'h18,
    8'h08,
    8'h04,
    8'h00,
    8'h00,
    8'h00,
    8'h10,
    8'h50,
    8'h2c,
    8'h38,
    8'h56,
    8'h10,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h18,
    8'h18,
    8'h18,
    8'hfe,
    8'h18,
    8'h18,
    8'h18,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h18,
    8'h18,
    8'h10,
    8'h0c,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h3c,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h18,
    8'h18,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h40,
    8'h60,
    8'h20,
    8'h30,
    8'h10,
    8'h10,
    8'h08,
    8'h08,
    8'h04,
    8'h04,
    8'h02,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h3c,
    8'h66,
    8'h42,
    8'he2,
    8'hda,
    8'hce,
    8'h42,
    8'h66,
    8'h3c,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h18,
    8'h1e,
    8'h12,
    8'h10,
    8'h10,
    8'h10,
    8'h10,
    8'h10,
    8'h7e,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h3c,
    8'h62,
    8'h60,
    8'h60,
    8'h20,
    8'h10,
    8'h08,
    8'h04,
    8'h7e,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h3e,
    8'h60,
    8'h60,
    8'h20,
    8'h3c,
    8'h40,
    8'h40,
    8'h60,
    8'h3e,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h30,
    8'h38,
    8'h28,
    8'h24,
    8'h26,
    8'h22,
    8'hff,
    8'h20,
    8'h20,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h7e,
    8'h06,
    8'h06,
    8'h06,
    8'h7e,
    8'h40,
    8'h40,
    8'h60,
    8'h3e,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h78,
    8'h0c,
    8'h06,
    8'h12,
    8'h6e,
    8'h42,
    8'h42,
    8'h46,
    8'h3c,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h7e,
    8'h40,
    8'h60,
    8'h20,
    8'h30,
    8'h10,
    8'h18,
    8'h08,
    8'h0c,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h3c,
    8'h46,
    8'h42,
    8'h6c,
    8'h38,
    8'h66,
    8'h42,
    8'h42,
    8'h3c,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h3c,
    8'h66,
    8'h42,
    8'h42,
    8'h66,
    8'h58,
    8'h40,
    8'h20,
    8'h1e,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h18,
    8'h18,
    8'h00,
    8'h00,
    8'h00,
    8'h18,
    8'h18,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h18,
    8'h18,
    8'h00,
    8'h00,
    8'h00,
    8'h18,
    8'h18,
    8'h10,
    8'h0c,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h20,
    8'h18,
    8'h0c,
    8'h06,
    8'h08,
    8'h30,
    8'h60,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h7e,
    8'h00,
    8'h7e,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h0c,
    8'h18,
    8'h20,
    8'h60,
    8'h30,
    8'h08,
    8'h04,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h0c,
    8'h38,
    8'h60,
    8'h60,
    8'h60,
    8'h18,
    8'h08,
    8'h00,
    8'h08,
    8'h08,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h38,
    8'h44,
    8'h82,
    8'h82,
    8'hbb,
    8'had,
    8'ha5,
    8'ha5,
    8'hf5,
    8'h29,
    8'h03,
    8'h02,
    8'h3c,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h18,
    8'h38,
    8'h2c,
    8'h24,
    8'h64,
    8'h46,
    8'h7e,
    8'hc2,
    8'h83,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h3e,
    8'h62,
    8'h42,
    8'h62,
    8'h3e,
    8'h42,
    8'h42,
    8'h42,
    8'h3e,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h78,
    8'h04,
    8'h02,
    8'h02,
    8'h02,
    8'h02,
    8'h02,
    8'h06,
    8'h7c,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h3e,
    8'h62,
    8'h42,
    8'hc2,
    8'hc2,
    8'hc2,
    8'h42,
    8'h62,
    8'h1e,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h7e,
    8'h06,
    8'h06,
    8'h06,
    8'h7e,
    8'h06,
    8'h06,
    8'h06,
    8'h7e,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h7e,
    8'h06,
    8'h06,
    8'h06,
    8'h7e,
    8'h06,
    8'h06,
    8'h06,
    8'h06,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h78,
    8'h06,
    8'h02,
    8'h02,
    8'h73,
    8'h42,
    8'h42,
    8'h46,
    8'h7c,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h42,
    8'h42,
    8'h42,
    8'h42,
    8'h7e,
    8'h42,
    8'h42,
    8'h42,
    8'h42,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h7e,
    8'h18,
    8'h18,
    8'h18,
    8'h18,
    8'h18,
    8'h18,
    8'h18,
    8'h7e,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h3e,
    8'h20,
    8'h20,
    8'h20,
    8'h20,
    8'h20,
    8'h20,
    8'h22,
    8'h1e,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h42,
    8'h22,
    8'h12,
    8'h0a,
    8'h0e,
    8'h1a,
    8'h32,
    8'h22,
    8'h42,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h04,
    8'h04,
    8'h04,
    8'h04,
    8'h04,
    8'h04,
    8'h04,
    8'h04,
    8'h7c,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h46,
    8'h66,
    8'he6,
    8'hfa,
    8'hda,
    8'hda,
    8'h83,
    8'h83,
    8'h83,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h46,
    8'h46,
    8'h4e,
    8'h4a,
    8'h5a,
    8'h52,
    8'h72,
    8'h62,
    8'h62,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h3c,
    8'h46,
    8'hc2,
    8'hc3,
    8'hc3,
    8'hc3,
    8'hc2,
    8'h46,
    8'h3c,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h3e,
    8'h62,
    8'h42,
    8'h42,
    8'h62,
    8'h1e,
    8'h02,
    8'h02,
    8'h02,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h3c,
    8'h46,
    8'hc2,
    8'hc3,
    8'hc3,
    8'hc3,
    8'hc2,
    8'h46,
    8'h3c,
    8'h18,
    8'hf0,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h3e,
    8'h66,
    8'h46,
    8'h66,
    8'h3e,
    8'h36,
    8'h26,
    8'h66,
    8'h46,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h7c,
    8'h06,
    8'h02,
    8'h06,
    8'h38,
    8'h60,
    8'h40,
    8'h40,
    8'h3e,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'hfe,
    8'h18,
    8'h18,
    8'h18,
    8'h18,
    8'h18,
    8'h18,
    8'h18,
    8'h18,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h42,
    8'h42,
    8'h42,
    8'h42,
    8'h42,
    8'h42,
    8'h42,
    8'h46,
    8'h3c,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h83,
    8'hc2,
    8'h42,
    8'h46,
    8'h64,
    8'h24,
    8'h2c,
    8'h38,
    8'h18,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h83,
    8'h83,
    8'h82,
    8'h92,
    8'hda,
    8'hda,
    8'h6e,
    8'h66,
    8'h66,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'hc2,
    8'h66,
    8'h2c,
    8'h18,
    8'h18,
    8'h38,
    8'h24,
    8'h66,
    8'hc3,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h83,
    8'h42,
    8'h66,
    8'h2c,
    8'h38,
    8'h18,
    8'h18,
    8'h18,
    8'h18,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h7e,
    8'h40,
    8'h20,
    8'h30,
    8'h18,
    8'h08,
    8'h04,
    8'h06,
    8'h7e,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h38,
    8'h08,
    8'h08,
    8'h08,
    8'h08,
    8'h08,
    8'h08,
    8'h08,
    8'h08,
    8'h08,
    8'h08,
    8'h08,
    8'h38,
    8'h00,
    8'h00,
    8'h00,
    8'h02,
    8'h04,
    8'h04,
    8'h08,
    8'h08,
    8'h10,
    8'h10,
    8'h30,
    8'h20,
    8'h60,
    8'h40,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h3c,
    8'h30,
    8'h30,
    8'h30,
    8'h30,
    8'h30,
    8'h30,
    8'h30,
    8'h30,
    8'h30,
    8'h30,
    8'h30,
    8'h3c,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h18,
    8'h38,
    8'h24,
    8'h46,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'hff,
    8'h00,
    8'h00,
    8'h00,
    8'h04,
    8'h08,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h3c,
    8'h60,
    8'h40,
    8'h7c,
    8'h42,
    8'h62,
    8'h5e,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h02,
    8'h02,
    8'h02,
    8'h3a,
    8'h46,
    8'h42,
    8'h42,
    8'h42,
    8'h42,
    8'h3e,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h78,
    8'h04,
    8'h06,
    8'h02,
    8'h06,
    8'h04,
    8'h7c,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h40,
    8'h40,
    8'h40,
    8'h7c,
    8'h46,
    8'h42,
    8'h42,
    8'h42,
    8'h66,
    8'h5c,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h3c,
    8'h46,
    8'h42,
    8'h7e,
    8'h02,
    8'h06,
    8'h7c,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'hf0,
    8'h18,
    8'h08,
    8'h08,
    8'h7e,
    8'h08,
    8'h08,
    8'h08,
    8'h08,
    8'h08,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'hfc,
    8'h66,
    8'h42,
    8'h66,
    8'h1a,
    8'h02,
    8'h7c,
    8'hc2,
    8'h42,
    8'h3c,
    8'h00,
    8'h00,
    8'h00,
    8'h02,
    8'h02,
    8'h02,
    8'h3a,
    8'h46,
    8'h42,
    8'h42,
    8'h42,
    8'h42,
    8'h42,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h18,
    8'h18,
    8'h00,
    8'h1e,
    8'h10,
    8'h10,
    8'h10,
    8'h10,
    8'h10,
    8'h7e,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h20,
    8'h30,
    8'h00,
    8'h3e,
    8'h20,
    8'h20,
    8'h20,
    8'h20,
    8'h20,
    8'h20,
    8'h20,
    8'h30,
    8'h1e,
    8'h00,
    8'h00,
    8'h00,
    8'h06,
    8'h06,
    8'h06,
    8'h46,
    8'h36,
    8'h1e,
    8'h0e,
    8'h16,
    8'h26,
    8'h46,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h1e,
    8'h10,
    8'h10,
    8'h10,
    8'h10,
    8'h10,
    8'h10,
    8'h10,
    8'h10,
    8'h7e,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h6e,
    8'hd2,
    8'hd2,
    8'hd2,
    8'hd2,
    8'hd2,
    8'hd2,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h3a,
    8'h46,
    8'h42,
    8'h42,
    8'h42,
    8'h42,
    8'h42,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h3c,
    8'h46,
    8'h42,
    8'hc2,
    8'h42,
    8'h46,
    8'h3c,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h3a,
    8'h46,
    8'h42,
    8'h42,
    8'h42,
    8'h42,
    8'h3e,
    8'h02,
    8'h02,
    8'h02,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h7c,
    8'h46,
    8'h42,
    8'h42,
    8'h42,
    8'h66,
    8'h5c,
    8'h40,
    8'h40,
    8'h40,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h76,
    8'h4e,
    8'hc6,
    8'h06,
    8'h06,
    8'h06,
    8'h06,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h7c,
    8'h04,
    8'h04,
    8'h3c,
    8'h60,
    8'h40,
    8'h3e,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h08,
    8'h08,
    8'h7f,
    8'h08,
    8'h08,
    8'h08,
    8'h08,
    8'h08,
    8'h78,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h42,
    8'h42,
    8'h42,
    8'h42,
    8'h42,
    8'h66,
    8'h5c,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'hc2,
    8'h42,
    8'h66,
    8'h24,
    8'h2c,
    8'h18,
    8'h18,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h83,
    8'h83,
    8'hda,
    8'h5a,
    8'h7a,
    8'h66,
    8'h66,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h46,
    8'h64,
    8'h38,
    8'h18,
    8'h38,
    8'h64,
    8'h46,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'hc2,
    8'h42,
    8'h66,
    8'h24,
    8'h2c,
    8'h38,
    8'h18,
    8'h18,
    8'h0c,
    8'h07,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h7e,
    8'h60,
    8'h30,
    8'h18,
    8'h08,
    8'h04,
    8'h7e,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h70,
    8'h18,
    8'h08,
    8'h08,
    8'h08,
    8'h0c,
    8'h0e,
    8'h08,
    8'h08,
    8'h08,
    8'h08,
    8'h18,
    8'h70,
    8'h00,
    8'h00,
    8'h10,
    8'h10,
    8'h10,
    8'h10,
    8'h10,
    8'h10,
    8'h10,
    8'h10,
    8'h10,
    8'h10,
    8'h10,
    8'h10,
    8'h10,
    8'h10,
    8'h00,
    8'h00,
    8'h00,
    8'h0c,
    8'h18,
    8'h10,
    8'h10,
    8'h10,
    8'h30,
    8'h70,
    8'h10,
    8'h10,
    8'h10,
    8'h10,
    8'h18,
    8'h0c,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h8e,
    8'hd2,
    8'h60,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00,
    8'h00
};

always @ (posedge clk)
    data <= rom_cell[addr];

endmodule

